//NOR gate using Structural modeling
module nor_gate_s(a,b,y);
input a,b;
output y;

nor(y,a,b);
                
endmodule