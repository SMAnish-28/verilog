//EX-OR gate using Structural modeling
module xor_gate_s(a,b,y);
input a,b;
output y;

xor(y,a,b);
                
endmodule