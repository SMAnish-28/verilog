//EX-NOR gate using Structural modeling
module xnor_gate_s(a,b,y);
input a,b;
output y;

xnor(y,a,b);
                
endmodule