//NAND gate using Structural modeling
module nand_gate_s(a,b,y);
input a,b;
output y;

nand(y,a,b);
                
endmodule