// NOT gate using structural modeling
module not_gate_s(a, y);
input a;
output y;

not(y, a); // syntax: gate_name(output, input)

endmodule